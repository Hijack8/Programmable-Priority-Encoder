module tothermo512(
  input [8:0] x,
  output [511:0] y
);
assign y[0] = ((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[1] = (((((((x[1]|x[2])|x[3])|x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[2] = ((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[3] = ((((((x[2]|x[3])|x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[4] = ((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[5] = (((((((x[1]&x[2])|x[3])|x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[6] = ((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[7] = (((((x[3]|x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[8] = ((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[9] = (((((((x[1]|x[2])&x[3])|x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[10] = ((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[11] = ((((((x[2]&x[3])|x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[12] = ((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[13] = (((((((x[1]&x[2])&x[3])|x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[14] = ((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[15] = ((((x[4]|x[5])|x[6])|x[7])|x[8]);
assign y[16] = ((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[17] = (((((((x[1]|x[2])|x[3])&x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[18] = ((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[19] = ((((((x[2]|x[3])&x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[20] = ((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[21] = (((((((x[1]&x[2])|x[3])&x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[22] = ((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[23] = (((((x[3]&x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[24] = ((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[25] = (((((((x[1]|x[2])&x[3])&x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[26] = ((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[27] = ((((((x[2]&x[3])&x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[28] = ((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[29] = (((((((x[1]&x[2])&x[3])&x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[30] = ((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])|x[6])|x[7])|x[8]);
assign y[31] = (((x[5]|x[6])|x[7])|x[8]);
assign y[32] = ((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[33] = (((((((x[1]|x[2])|x[3])|x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[34] = ((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[35] = ((((((x[2]|x[3])|x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[36] = ((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[37] = (((((((x[1]&x[2])|x[3])|x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[38] = ((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[39] = (((((x[3]|x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[40] = ((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[41] = (((((((x[1]|x[2])&x[3])|x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[42] = ((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[43] = ((((((x[2]&x[3])|x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[44] = ((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[45] = (((((((x[1]&x[2])&x[3])|x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[46] = ((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[47] = ((((x[4]&x[5])|x[6])|x[7])|x[8]);
assign y[48] = ((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[49] = (((((((x[1]|x[2])|x[3])&x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[50] = ((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[51] = ((((((x[2]|x[3])&x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[52] = ((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[53] = (((((((x[1]&x[2])|x[3])&x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[54] = ((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[55] = (((((x[3]&x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[56] = ((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[57] = (((((((x[1]|x[2])&x[3])&x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[58] = ((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[59] = ((((((x[2]&x[3])&x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[60] = ((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[61] = (((((((x[1]&x[2])&x[3])&x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[62] = ((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])|x[6])|x[7])|x[8]);
assign y[63] = ((x[6]|x[7])|x[8]);
assign y[64] = ((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[65] = (((((((x[1]|x[2])|x[3])|x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[66] = ((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[67] = ((((((x[2]|x[3])|x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[68] = ((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[69] = (((((((x[1]&x[2])|x[3])|x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[70] = ((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[71] = (((((x[3]|x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[72] = ((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[73] = (((((((x[1]|x[2])&x[3])|x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[74] = ((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[75] = ((((((x[2]&x[3])|x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[76] = ((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[77] = (((((((x[1]&x[2])&x[3])|x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[78] = ((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[79] = ((((x[4]|x[5])&x[6])|x[7])|x[8]);
assign y[80] = ((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[81] = (((((((x[1]|x[2])|x[3])&x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[82] = ((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[83] = ((((((x[2]|x[3])&x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[84] = ((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[85] = (((((((x[1]&x[2])|x[3])&x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[86] = ((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[87] = (((((x[3]&x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[88] = ((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[89] = (((((((x[1]|x[2])&x[3])&x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[90] = ((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[91] = ((((((x[2]&x[3])&x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[92] = ((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[93] = (((((((x[1]&x[2])&x[3])&x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[94] = ((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])&x[6])|x[7])|x[8]);
assign y[95] = (((x[5]&x[6])|x[7])|x[8]);
assign y[96] = ((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[97] = (((((((x[1]|x[2])|x[3])|x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[98] = ((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[99] = ((((((x[2]|x[3])|x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[100] = ((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[101] = (((((((x[1]&x[2])|x[3])|x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[102] = ((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[103] = (((((x[3]|x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[104] = ((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[105] = (((((((x[1]|x[2])&x[3])|x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[106] = ((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[107] = ((((((x[2]&x[3])|x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[108] = ((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[109] = (((((((x[1]&x[2])&x[3])|x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[110] = ((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[111] = ((((x[4]&x[5])&x[6])|x[7])|x[8]);
assign y[112] = ((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[113] = (((((((x[1]|x[2])|x[3])&x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[114] = ((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[115] = ((((((x[2]|x[3])&x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[116] = ((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[117] = (((((((x[1]&x[2])|x[3])&x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[118] = ((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[119] = (((((x[3]&x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[120] = ((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[121] = (((((((x[1]|x[2])&x[3])&x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[122] = ((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[123] = ((((((x[2]&x[3])&x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[124] = ((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[125] = (((((((x[1]&x[2])&x[3])&x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[126] = ((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])&x[6])|x[7])|x[8]);
assign y[127] = (x[7]|x[8]);
assign y[128] = ((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[129] = (((((((x[1]|x[2])|x[3])|x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[130] = ((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[131] = ((((((x[2]|x[3])|x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[132] = ((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[133] = (((((((x[1]&x[2])|x[3])|x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[134] = ((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[135] = (((((x[3]|x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[136] = ((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[137] = (((((((x[1]|x[2])&x[3])|x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[138] = ((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[139] = ((((((x[2]&x[3])|x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[140] = ((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[141] = (((((((x[1]&x[2])&x[3])|x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[142] = ((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[143] = ((((x[4]|x[5])|x[6])&x[7])|x[8]);
assign y[144] = ((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[145] = (((((((x[1]|x[2])|x[3])&x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[146] = ((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[147] = ((((((x[2]|x[3])&x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[148] = ((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[149] = (((((((x[1]&x[2])|x[3])&x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[150] = ((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[151] = (((((x[3]&x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[152] = ((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[153] = (((((((x[1]|x[2])&x[3])&x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[154] = ((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[155] = ((((((x[2]&x[3])&x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[156] = ((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[157] = (((((((x[1]&x[2])&x[3])&x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[158] = ((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])|x[6])&x[7])|x[8]);
assign y[159] = (((x[5]|x[6])&x[7])|x[8]);
assign y[160] = ((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[161] = (((((((x[1]|x[2])|x[3])|x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[162] = ((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[163] = ((((((x[2]|x[3])|x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[164] = ((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[165] = (((((((x[1]&x[2])|x[3])|x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[166] = ((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[167] = (((((x[3]|x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[168] = ((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[169] = (((((((x[1]|x[2])&x[3])|x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[170] = ((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[171] = ((((((x[2]&x[3])|x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[172] = ((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[173] = (((((((x[1]&x[2])&x[3])|x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[174] = ((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[175] = ((((x[4]&x[5])|x[6])&x[7])|x[8]);
assign y[176] = ((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[177] = (((((((x[1]|x[2])|x[3])&x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[178] = ((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[179] = ((((((x[2]|x[3])&x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[180] = ((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[181] = (((((((x[1]&x[2])|x[3])&x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[182] = ((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[183] = (((((x[3]&x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[184] = ((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[185] = (((((((x[1]|x[2])&x[3])&x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[186] = ((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[187] = ((((((x[2]&x[3])&x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[188] = ((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[189] = (((((((x[1]&x[2])&x[3])&x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[190] = ((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])|x[6])&x[7])|x[8]);
assign y[191] = ((x[6]&x[7])|x[8]);
assign y[192] = ((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[193] = (((((((x[1]|x[2])|x[3])|x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[194] = ((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[195] = ((((((x[2]|x[3])|x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[196] = ((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[197] = (((((((x[1]&x[2])|x[3])|x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[198] = ((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[199] = (((((x[3]|x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[200] = ((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[201] = (((((((x[1]|x[2])&x[3])|x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[202] = ((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[203] = ((((((x[2]&x[3])|x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[204] = ((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[205] = (((((((x[1]&x[2])&x[3])|x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[206] = ((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[207] = ((((x[4]|x[5])&x[6])&x[7])|x[8]);
assign y[208] = ((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[209] = (((((((x[1]|x[2])|x[3])&x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[210] = ((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[211] = ((((((x[2]|x[3])&x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[212] = ((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[213] = (((((((x[1]&x[2])|x[3])&x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[214] = ((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[215] = (((((x[3]&x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[216] = ((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[217] = (((((((x[1]|x[2])&x[3])&x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[218] = ((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[219] = ((((((x[2]&x[3])&x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[220] = ((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[221] = (((((((x[1]&x[2])&x[3])&x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[222] = ((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])&x[6])&x[7])|x[8]);
assign y[223] = (((x[5]&x[6])&x[7])|x[8]);
assign y[224] = ((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[225] = (((((((x[1]|x[2])|x[3])|x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[226] = ((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[227] = ((((((x[2]|x[3])|x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[228] = ((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[229] = (((((((x[1]&x[2])|x[3])|x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[230] = ((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[231] = (((((x[3]|x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[232] = ((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[233] = (((((((x[1]|x[2])&x[3])|x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[234] = ((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[235] = ((((((x[2]&x[3])|x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[236] = ((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[237] = (((((((x[1]&x[2])&x[3])|x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[238] = ((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[239] = ((((x[4]&x[5])&x[6])&x[7])|x[8]);
assign y[240] = ((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[241] = (((((((x[1]|x[2])|x[3])&x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[242] = ((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[243] = ((((((x[2]|x[3])&x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[244] = ((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[245] = (((((((x[1]&x[2])|x[3])&x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[246] = ((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[247] = (((((x[3]&x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[248] = ((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[249] = (((((((x[1]|x[2])&x[3])&x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[250] = ((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[251] = ((((((x[2]&x[3])&x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[252] = ((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[253] = (((((((x[1]&x[2])&x[3])&x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[254] = ((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])&x[6])&x[7])|x[8]);
assign y[255] = x[8];
assign y[256] = ((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[257] = (((((((x[1]|x[2])|x[3])|x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[258] = ((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[259] = ((((((x[2]|x[3])|x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[260] = ((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[261] = (((((((x[1]&x[2])|x[3])|x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[262] = ((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[263] = (((((x[3]|x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[264] = ((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[265] = (((((((x[1]|x[2])&x[3])|x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[266] = ((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[267] = ((((((x[2]&x[3])|x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[268] = ((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[269] = (((((((x[1]&x[2])&x[3])|x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[270] = ((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[271] = ((((x[4]|x[5])|x[6])|x[7])&x[8]);
assign y[272] = ((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[273] = (((((((x[1]|x[2])|x[3])&x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[274] = ((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[275] = ((((((x[2]|x[3])&x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[276] = ((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[277] = (((((((x[1]&x[2])|x[3])&x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[278] = ((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[279] = (((((x[3]&x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[280] = ((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[281] = (((((((x[1]|x[2])&x[3])&x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[282] = ((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[283] = ((((((x[2]&x[3])&x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[284] = ((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[285] = (((((((x[1]&x[2])&x[3])&x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[286] = ((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])|x[6])|x[7])&x[8]);
assign y[287] = (((x[5]|x[6])|x[7])&x[8]);
assign y[288] = ((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[289] = (((((((x[1]|x[2])|x[3])|x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[290] = ((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[291] = ((((((x[2]|x[3])|x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[292] = ((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[293] = (((((((x[1]&x[2])|x[3])|x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[294] = ((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[295] = (((((x[3]|x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[296] = ((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[297] = (((((((x[1]|x[2])&x[3])|x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[298] = ((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[299] = ((((((x[2]&x[3])|x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[300] = ((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[301] = (((((((x[1]&x[2])&x[3])|x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[302] = ((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[303] = ((((x[4]&x[5])|x[6])|x[7])&x[8]);
assign y[304] = ((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[305] = (((((((x[1]|x[2])|x[3])&x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[306] = ((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[307] = ((((((x[2]|x[3])&x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[308] = ((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[309] = (((((((x[1]&x[2])|x[3])&x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[310] = ((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[311] = (((((x[3]&x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[312] = ((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[313] = (((((((x[1]|x[2])&x[3])&x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[314] = ((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[315] = ((((((x[2]&x[3])&x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[316] = ((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[317] = (((((((x[1]&x[2])&x[3])&x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[318] = ((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])|x[6])|x[7])&x[8]);
assign y[319] = ((x[6]|x[7])&x[8]);
assign y[320] = ((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[321] = (((((((x[1]|x[2])|x[3])|x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[322] = ((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[323] = ((((((x[2]|x[3])|x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[324] = ((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[325] = (((((((x[1]&x[2])|x[3])|x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[326] = ((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[327] = (((((x[3]|x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[328] = ((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[329] = (((((((x[1]|x[2])&x[3])|x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[330] = ((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[331] = ((((((x[2]&x[3])|x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[332] = ((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[333] = (((((((x[1]&x[2])&x[3])|x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[334] = ((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[335] = ((((x[4]|x[5])&x[6])|x[7])&x[8]);
assign y[336] = ((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[337] = (((((((x[1]|x[2])|x[3])&x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[338] = ((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[339] = ((((((x[2]|x[3])&x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[340] = ((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[341] = (((((((x[1]&x[2])|x[3])&x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[342] = ((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[343] = (((((x[3]&x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[344] = ((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[345] = (((((((x[1]|x[2])&x[3])&x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[346] = ((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[347] = ((((((x[2]&x[3])&x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[348] = ((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[349] = (((((((x[1]&x[2])&x[3])&x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[350] = ((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])&x[6])|x[7])&x[8]);
assign y[351] = (((x[5]&x[6])|x[7])&x[8]);
assign y[352] = ((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[353] = (((((((x[1]|x[2])|x[3])|x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[354] = ((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[355] = ((((((x[2]|x[3])|x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[356] = ((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[357] = (((((((x[1]&x[2])|x[3])|x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[358] = ((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[359] = (((((x[3]|x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[360] = ((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[361] = (((((((x[1]|x[2])&x[3])|x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[362] = ((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[363] = ((((((x[2]&x[3])|x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[364] = ((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[365] = (((((((x[1]&x[2])&x[3])|x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[366] = ((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[367] = ((((x[4]&x[5])&x[6])|x[7])&x[8]);
assign y[368] = ((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[369] = (((((((x[1]|x[2])|x[3])&x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[370] = ((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[371] = ((((((x[2]|x[3])&x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[372] = ((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[373] = (((((((x[1]&x[2])|x[3])&x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[374] = ((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[375] = (((((x[3]&x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[376] = ((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[377] = (((((((x[1]|x[2])&x[3])&x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[378] = ((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[379] = ((((((x[2]&x[3])&x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[380] = ((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[381] = (((((((x[1]&x[2])&x[3])&x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[382] = ((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])&x[6])|x[7])&x[8]);
assign y[383] = (x[7]&x[8]);
assign y[384] = ((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[385] = (((((((x[1]|x[2])|x[3])|x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[386] = ((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[387] = ((((((x[2]|x[3])|x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[388] = ((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[389] = (((((((x[1]&x[2])|x[3])|x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[390] = ((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[391] = (((((x[3]|x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[392] = ((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[393] = (((((((x[1]|x[2])&x[3])|x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[394] = ((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[395] = ((((((x[2]&x[3])|x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[396] = ((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[397] = (((((((x[1]&x[2])&x[3])|x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[398] = ((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[399] = ((((x[4]|x[5])|x[6])&x[7])&x[8]);
assign y[400] = ((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[401] = (((((((x[1]|x[2])|x[3])&x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[402] = ((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[403] = ((((((x[2]|x[3])&x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[404] = ((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[405] = (((((((x[1]&x[2])|x[3])&x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[406] = ((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[407] = (((((x[3]&x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[408] = ((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[409] = (((((((x[1]|x[2])&x[3])&x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[410] = ((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[411] = ((((((x[2]&x[3])&x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[412] = ((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[413] = (((((((x[1]&x[2])&x[3])&x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[414] = ((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])|x[6])&x[7])&x[8]);
assign y[415] = (((x[5]|x[6])&x[7])&x[8]);
assign y[416] = ((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[417] = (((((((x[1]|x[2])|x[3])|x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[418] = ((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[419] = ((((((x[2]|x[3])|x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[420] = ((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[421] = (((((((x[1]&x[2])|x[3])|x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[422] = ((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[423] = (((((x[3]|x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[424] = ((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[425] = (((((((x[1]|x[2])&x[3])|x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[426] = ((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[427] = ((((((x[2]&x[3])|x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[428] = ((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[429] = (((((((x[1]&x[2])&x[3])|x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[430] = ((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[431] = ((((x[4]&x[5])|x[6])&x[7])&x[8]);
assign y[432] = ((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[433] = (((((((x[1]|x[2])|x[3])&x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[434] = ((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[435] = ((((((x[2]|x[3])&x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[436] = ((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[437] = (((((((x[1]&x[2])|x[3])&x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[438] = ((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[439] = (((((x[3]&x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[440] = ((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[441] = (((((((x[1]|x[2])&x[3])&x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[442] = ((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[443] = ((((((x[2]&x[3])&x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[444] = ((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[445] = (((((((x[1]&x[2])&x[3])&x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[446] = ((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])|x[6])&x[7])&x[8]);
assign y[447] = ((x[6]&x[7])&x[8]);
assign y[448] = ((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[449] = (((((((x[1]|x[2])|x[3])|x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[450] = ((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[451] = ((((((x[2]|x[3])|x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[452] = ((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[453] = (((((((x[1]&x[2])|x[3])|x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[454] = ((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[455] = (((((x[3]|x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[456] = ((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[457] = (((((((x[1]|x[2])&x[3])|x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[458] = ((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[459] = ((((((x[2]&x[3])|x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[460] = ((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[461] = (((((((x[1]&x[2])&x[3])|x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[462] = ((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[463] = ((((x[4]|x[5])&x[6])&x[7])&x[8]);
assign y[464] = ((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[465] = (((((((x[1]|x[2])|x[3])&x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[466] = ((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[467] = ((((((x[2]|x[3])&x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[468] = ((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[469] = (((((((x[1]&x[2])|x[3])&x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[470] = ((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[471] = (((((x[3]&x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[472] = ((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[473] = (((((((x[1]|x[2])&x[3])&x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[474] = ((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[475] = ((((((x[2]&x[3])&x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[476] = ((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[477] = (((((((x[1]&x[2])&x[3])&x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[478] = ((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])&x[6])&x[7])&x[8]);
assign y[479] = (((x[5]&x[6])&x[7])&x[8]);
assign y[480] = ((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[481] = (((((((x[1]|x[2])|x[3])|x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[482] = ((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[483] = ((((((x[2]|x[3])|x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[484] = ((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[485] = (((((((x[1]&x[2])|x[3])|x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[486] = ((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[487] = (((((x[3]|x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[488] = ((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[489] = (((((((x[1]|x[2])&x[3])|x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[490] = ((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[491] = ((((((x[2]&x[3])|x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[492] = ((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[493] = (((((((x[1]&x[2])&x[3])|x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[494] = ((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[495] = ((((x[4]&x[5])&x[6])&x[7])&x[8]);
assign y[496] = ((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[497] = (((((((x[1]|x[2])|x[3])&x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[498] = ((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[499] = ((((((x[2]|x[3])&x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[500] = ((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[501] = (((((((x[1]&x[2])|x[3])&x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[502] = ((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[503] = (((((x[3]&x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[504] = ((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[505] = (((((((x[1]|x[2])&x[3])&x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[506] = ((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[507] = ((((((x[2]&x[3])&x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[508] = ((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[509] = (((((((x[1]&x[2])&x[3])&x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[510] = ((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])&x[6])&x[7])&x[8]);
assign y[511] = 0;
endmodule 
