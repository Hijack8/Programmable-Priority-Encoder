
module tothermo1024(
  input [9:0] x,
  output [1023:0] y
);

assign y[0] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[1] = ((((((((x[1]|x[2])|x[3])|x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[2] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[3] = (((((((x[2]|x[3])|x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[4] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[5] = ((((((((x[1]&x[2])|x[3])|x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[6] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[7] = ((((((x[3]|x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[8] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[9] = ((((((((x[1]|x[2])&x[3])|x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[10] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[11] = (((((((x[2]&x[3])|x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[12] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[13] = ((((((((x[1]&x[2])&x[3])|x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[14] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[15] = (((((x[4]|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[16] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[17] = ((((((((x[1]|x[2])|x[3])&x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[18] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[19] = (((((((x[2]|x[3])&x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[20] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[21] = ((((((((x[1]&x[2])|x[3])&x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[22] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[23] = ((((((x[3]&x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[24] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[25] = ((((((((x[1]|x[2])&x[3])&x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[26] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[27] = (((((((x[2]&x[3])&x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[28] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[29] = ((((((((x[1]&x[2])&x[3])&x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[30] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[31] = ((((x[5]|x[6])|x[7])|x[8])|x[9]);
assign y[32] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[33] = ((((((((x[1]|x[2])|x[3])|x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[34] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[35] = (((((((x[2]|x[3])|x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[36] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[37] = ((((((((x[1]&x[2])|x[3])|x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[38] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[39] = ((((((x[3]|x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[40] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[41] = ((((((((x[1]|x[2])&x[3])|x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[42] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[43] = (((((((x[2]&x[3])|x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[44] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[45] = ((((((((x[1]&x[2])&x[3])|x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[46] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[47] = (((((x[4]&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[48] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[49] = ((((((((x[1]|x[2])|x[3])&x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[50] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[51] = (((((((x[2]|x[3])&x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[52] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[53] = ((((((((x[1]&x[2])|x[3])&x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[54] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[55] = ((((((x[3]&x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[56] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[57] = ((((((((x[1]|x[2])&x[3])&x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[58] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[59] = (((((((x[2]&x[3])&x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[60] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[61] = ((((((((x[1]&x[2])&x[3])&x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[62] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])|x[6])|x[7])|x[8])|x[9]);
assign y[63] = (((x[6]|x[7])|x[8])|x[9]);
assign y[64] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[65] = ((((((((x[1]|x[2])|x[3])|x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[66] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[67] = (((((((x[2]|x[3])|x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[68] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[69] = ((((((((x[1]&x[2])|x[3])|x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[70] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[71] = ((((((x[3]|x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[72] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[73] = ((((((((x[1]|x[2])&x[3])|x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[74] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[75] = (((((((x[2]&x[3])|x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[76] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[77] = ((((((((x[1]&x[2])&x[3])|x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[78] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[79] = (((((x[4]|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[80] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[81] = ((((((((x[1]|x[2])|x[3])&x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[82] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[83] = (((((((x[2]|x[3])&x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[84] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[85] = ((((((((x[1]&x[2])|x[3])&x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[86] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[87] = ((((((x[3]&x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[88] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[89] = ((((((((x[1]|x[2])&x[3])&x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[90] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[91] = (((((((x[2]&x[3])&x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[92] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[93] = ((((((((x[1]&x[2])&x[3])&x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[94] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[95] = ((((x[5]&x[6])|x[7])|x[8])|x[9]);
assign y[96] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[97] = ((((((((x[1]|x[2])|x[3])|x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[98] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[99] = (((((((x[2]|x[3])|x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[100] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[101] = ((((((((x[1]&x[2])|x[3])|x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[102] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[103] = ((((((x[3]|x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[104] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[105] = ((((((((x[1]|x[2])&x[3])|x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[106] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[107] = (((((((x[2]&x[3])|x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[108] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[109] = ((((((((x[1]&x[2])&x[3])|x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[110] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[111] = (((((x[4]&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[112] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[113] = ((((((((x[1]|x[2])|x[3])&x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[114] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[115] = (((((((x[2]|x[3])&x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[116] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[117] = ((((((((x[1]&x[2])|x[3])&x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[118] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[119] = ((((((x[3]&x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[120] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[121] = ((((((((x[1]|x[2])&x[3])&x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[122] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[123] = (((((((x[2]&x[3])&x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[124] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[125] = ((((((((x[1]&x[2])&x[3])&x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[126] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])&x[6])|x[7])|x[8])|x[9]);
assign y[127] = ((x[7]|x[8])|x[9]);
assign y[128] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[129] = ((((((((x[1]|x[2])|x[3])|x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[130] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[131] = (((((((x[2]|x[3])|x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[132] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[133] = ((((((((x[1]&x[2])|x[3])|x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[134] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[135] = ((((((x[3]|x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[136] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[137] = ((((((((x[1]|x[2])&x[3])|x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[138] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[139] = (((((((x[2]&x[3])|x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[140] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[141] = ((((((((x[1]&x[2])&x[3])|x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[142] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[143] = (((((x[4]|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[144] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[145] = ((((((((x[1]|x[2])|x[3])&x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[146] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[147] = (((((((x[2]|x[3])&x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[148] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[149] = ((((((((x[1]&x[2])|x[3])&x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[150] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[151] = ((((((x[3]&x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[152] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[153] = ((((((((x[1]|x[2])&x[3])&x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[154] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[155] = (((((((x[2]&x[3])&x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[156] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[157] = ((((((((x[1]&x[2])&x[3])&x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[158] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[159] = ((((x[5]|x[6])&x[7])|x[8])|x[9]);
assign y[160] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[161] = ((((((((x[1]|x[2])|x[3])|x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[162] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[163] = (((((((x[2]|x[3])|x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[164] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[165] = ((((((((x[1]&x[2])|x[3])|x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[166] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[167] = ((((((x[3]|x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[168] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[169] = ((((((((x[1]|x[2])&x[3])|x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[170] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[171] = (((((((x[2]&x[3])|x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[172] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[173] = ((((((((x[1]&x[2])&x[3])|x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[174] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[175] = (((((x[4]&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[176] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[177] = ((((((((x[1]|x[2])|x[3])&x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[178] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[179] = (((((((x[2]|x[3])&x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[180] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[181] = ((((((((x[1]&x[2])|x[3])&x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[182] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[183] = ((((((x[3]&x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[184] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[185] = ((((((((x[1]|x[2])&x[3])&x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[186] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[187] = (((((((x[2]&x[3])&x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[188] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[189] = ((((((((x[1]&x[2])&x[3])&x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[190] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])|x[6])&x[7])|x[8])|x[9]);
assign y[191] = (((x[6]&x[7])|x[8])|x[9]);
assign y[192] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[193] = ((((((((x[1]|x[2])|x[3])|x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[194] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[195] = (((((((x[2]|x[3])|x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[196] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[197] = ((((((((x[1]&x[2])|x[3])|x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[198] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[199] = ((((((x[3]|x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[200] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[201] = ((((((((x[1]|x[2])&x[3])|x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[202] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[203] = (((((((x[2]&x[3])|x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[204] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[205] = ((((((((x[1]&x[2])&x[3])|x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[206] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[207] = (((((x[4]|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[208] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[209] = ((((((((x[1]|x[2])|x[3])&x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[210] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[211] = (((((((x[2]|x[3])&x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[212] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[213] = ((((((((x[1]&x[2])|x[3])&x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[214] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[215] = ((((((x[3]&x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[216] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[217] = ((((((((x[1]|x[2])&x[3])&x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[218] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[219] = (((((((x[2]&x[3])&x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[220] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[221] = ((((((((x[1]&x[2])&x[3])&x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[222] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[223] = ((((x[5]&x[6])&x[7])|x[8])|x[9]);
assign y[224] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[225] = ((((((((x[1]|x[2])|x[3])|x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[226] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[227] = (((((((x[2]|x[3])|x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[228] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[229] = ((((((((x[1]&x[2])|x[3])|x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[230] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[231] = ((((((x[3]|x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[232] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[233] = ((((((((x[1]|x[2])&x[3])|x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[234] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[235] = (((((((x[2]&x[3])|x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[236] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[237] = ((((((((x[1]&x[2])&x[3])|x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[238] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[239] = (((((x[4]&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[240] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[241] = ((((((((x[1]|x[2])|x[3])&x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[242] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[243] = (((((((x[2]|x[3])&x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[244] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[245] = ((((((((x[1]&x[2])|x[3])&x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[246] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[247] = ((((((x[3]&x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[248] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[249] = ((((((((x[1]|x[2])&x[3])&x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[250] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[251] = (((((((x[2]&x[3])&x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[252] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[253] = ((((((((x[1]&x[2])&x[3])&x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[254] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])&x[6])&x[7])|x[8])|x[9]);
assign y[255] = (x[8]|x[9]);
assign y[256] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[257] = ((((((((x[1]|x[2])|x[3])|x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[258] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[259] = (((((((x[2]|x[3])|x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[260] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[261] = ((((((((x[1]&x[2])|x[3])|x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[262] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[263] = ((((((x[3]|x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[264] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[265] = ((((((((x[1]|x[2])&x[3])|x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[266] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[267] = (((((((x[2]&x[3])|x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[268] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[269] = ((((((((x[1]&x[2])&x[3])|x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[270] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[271] = (((((x[4]|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[272] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[273] = ((((((((x[1]|x[2])|x[3])&x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[274] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[275] = (((((((x[2]|x[3])&x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[276] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[277] = ((((((((x[1]&x[2])|x[3])&x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[278] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[279] = ((((((x[3]&x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[280] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[281] = ((((((((x[1]|x[2])&x[3])&x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[282] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[283] = (((((((x[2]&x[3])&x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[284] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[285] = ((((((((x[1]&x[2])&x[3])&x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[286] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[287] = ((((x[5]|x[6])|x[7])&x[8])|x[9]);
assign y[288] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[289] = ((((((((x[1]|x[2])|x[3])|x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[290] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[291] = (((((((x[2]|x[3])|x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[292] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[293] = ((((((((x[1]&x[2])|x[3])|x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[294] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[295] = ((((((x[3]|x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[296] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[297] = ((((((((x[1]|x[2])&x[3])|x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[298] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[299] = (((((((x[2]&x[3])|x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[300] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[301] = ((((((((x[1]&x[2])&x[3])|x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[302] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[303] = (((((x[4]&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[304] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[305] = ((((((((x[1]|x[2])|x[3])&x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[306] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[307] = (((((((x[2]|x[3])&x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[308] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[309] = ((((((((x[1]&x[2])|x[3])&x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[310] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[311] = ((((((x[3]&x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[312] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[313] = ((((((((x[1]|x[2])&x[3])&x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[314] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[315] = (((((((x[2]&x[3])&x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[316] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[317] = ((((((((x[1]&x[2])&x[3])&x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[318] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])|x[6])|x[7])&x[8])|x[9]);
assign y[319] = (((x[6]|x[7])&x[8])|x[9]);
assign y[320] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[321] = ((((((((x[1]|x[2])|x[3])|x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[322] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[323] = (((((((x[2]|x[3])|x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[324] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[325] = ((((((((x[1]&x[2])|x[3])|x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[326] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[327] = ((((((x[3]|x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[328] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[329] = ((((((((x[1]|x[2])&x[3])|x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[330] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[331] = (((((((x[2]&x[3])|x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[332] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[333] = ((((((((x[1]&x[2])&x[3])|x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[334] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[335] = (((((x[4]|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[336] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[337] = ((((((((x[1]|x[2])|x[3])&x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[338] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[339] = (((((((x[2]|x[3])&x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[340] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[341] = ((((((((x[1]&x[2])|x[3])&x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[342] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[343] = ((((((x[3]&x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[344] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[345] = ((((((((x[1]|x[2])&x[3])&x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[346] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[347] = (((((((x[2]&x[3])&x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[348] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[349] = ((((((((x[1]&x[2])&x[3])&x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[350] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[351] = ((((x[5]&x[6])|x[7])&x[8])|x[9]);
assign y[352] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[353] = ((((((((x[1]|x[2])|x[3])|x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[354] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[355] = (((((((x[2]|x[3])|x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[356] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[357] = ((((((((x[1]&x[2])|x[3])|x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[358] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[359] = ((((((x[3]|x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[360] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[361] = ((((((((x[1]|x[2])&x[3])|x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[362] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[363] = (((((((x[2]&x[3])|x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[364] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[365] = ((((((((x[1]&x[2])&x[3])|x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[366] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[367] = (((((x[4]&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[368] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[369] = ((((((((x[1]|x[2])|x[3])&x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[370] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[371] = (((((((x[2]|x[3])&x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[372] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[373] = ((((((((x[1]&x[2])|x[3])&x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[374] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[375] = ((((((x[3]&x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[376] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[377] = ((((((((x[1]|x[2])&x[3])&x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[378] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[379] = (((((((x[2]&x[3])&x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[380] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[381] = ((((((((x[1]&x[2])&x[3])&x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[382] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])&x[6])|x[7])&x[8])|x[9]);
assign y[383] = ((x[7]&x[8])|x[9]);
assign y[384] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[385] = ((((((((x[1]|x[2])|x[3])|x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[386] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[387] = (((((((x[2]|x[3])|x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[388] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[389] = ((((((((x[1]&x[2])|x[3])|x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[390] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[391] = ((((((x[3]|x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[392] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[393] = ((((((((x[1]|x[2])&x[3])|x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[394] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[395] = (((((((x[2]&x[3])|x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[396] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[397] = ((((((((x[1]&x[2])&x[3])|x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[398] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[399] = (((((x[4]|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[400] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[401] = ((((((((x[1]|x[2])|x[3])&x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[402] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[403] = (((((((x[2]|x[3])&x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[404] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[405] = ((((((((x[1]&x[2])|x[3])&x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[406] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[407] = ((((((x[3]&x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[408] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[409] = ((((((((x[1]|x[2])&x[3])&x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[410] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[411] = (((((((x[2]&x[3])&x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[412] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[413] = ((((((((x[1]&x[2])&x[3])&x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[414] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[415] = ((((x[5]|x[6])&x[7])&x[8])|x[9]);
assign y[416] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[417] = ((((((((x[1]|x[2])|x[3])|x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[418] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[419] = (((((((x[2]|x[3])|x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[420] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[421] = ((((((((x[1]&x[2])|x[3])|x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[422] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[423] = ((((((x[3]|x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[424] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[425] = ((((((((x[1]|x[2])&x[3])|x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[426] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[427] = (((((((x[2]&x[3])|x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[428] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[429] = ((((((((x[1]&x[2])&x[3])|x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[430] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[431] = (((((x[4]&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[432] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[433] = ((((((((x[1]|x[2])|x[3])&x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[434] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[435] = (((((((x[2]|x[3])&x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[436] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[437] = ((((((((x[1]&x[2])|x[3])&x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[438] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[439] = ((((((x[3]&x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[440] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[441] = ((((((((x[1]|x[2])&x[3])&x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[442] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[443] = (((((((x[2]&x[3])&x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[444] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[445] = ((((((((x[1]&x[2])&x[3])&x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[446] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])|x[6])&x[7])&x[8])|x[9]);
assign y[447] = (((x[6]&x[7])&x[8])|x[9]);
assign y[448] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[449] = ((((((((x[1]|x[2])|x[3])|x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[450] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[451] = (((((((x[2]|x[3])|x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[452] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[453] = ((((((((x[1]&x[2])|x[3])|x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[454] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[455] = ((((((x[3]|x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[456] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[457] = ((((((((x[1]|x[2])&x[3])|x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[458] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[459] = (((((((x[2]&x[3])|x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[460] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[461] = ((((((((x[1]&x[2])&x[3])|x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[462] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[463] = (((((x[4]|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[464] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[465] = ((((((((x[1]|x[2])|x[3])&x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[466] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[467] = (((((((x[2]|x[3])&x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[468] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[469] = ((((((((x[1]&x[2])|x[3])&x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[470] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[471] = ((((((x[3]&x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[472] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[473] = ((((((((x[1]|x[2])&x[3])&x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[474] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[475] = (((((((x[2]&x[3])&x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[476] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[477] = ((((((((x[1]&x[2])&x[3])&x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[478] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[479] = ((((x[5]&x[6])&x[7])&x[8])|x[9]);
assign y[480] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[481] = ((((((((x[1]|x[2])|x[3])|x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[482] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[483] = (((((((x[2]|x[3])|x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[484] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[485] = ((((((((x[1]&x[2])|x[3])|x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[486] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[487] = ((((((x[3]|x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[488] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[489] = ((((((((x[1]|x[2])&x[3])|x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[490] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[491] = (((((((x[2]&x[3])|x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[492] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[493] = ((((((((x[1]&x[2])&x[3])|x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[494] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[495] = (((((x[4]&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[496] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[497] = ((((((((x[1]|x[2])|x[3])&x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[498] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[499] = (((((((x[2]|x[3])&x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[500] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[501] = ((((((((x[1]&x[2])|x[3])&x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[502] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[503] = ((((((x[3]&x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[504] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[505] = ((((((((x[1]|x[2])&x[3])&x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[506] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[507] = (((((((x[2]&x[3])&x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[508] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[509] = ((((((((x[1]&x[2])&x[3])&x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[510] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])&x[6])&x[7])&x[8])|x[9]);
assign y[511] = x[9];
assign y[512] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[513] = ((((((((x[1]|x[2])|x[3])|x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[514] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[515] = (((((((x[2]|x[3])|x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[516] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[517] = ((((((((x[1]&x[2])|x[3])|x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[518] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[519] = ((((((x[3]|x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[520] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[521] = ((((((((x[1]|x[2])&x[3])|x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[522] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[523] = (((((((x[2]&x[3])|x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[524] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[525] = ((((((((x[1]&x[2])&x[3])|x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[526] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[527] = (((((x[4]|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[528] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[529] = ((((((((x[1]|x[2])|x[3])&x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[530] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[531] = (((((((x[2]|x[3])&x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[532] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[533] = ((((((((x[1]&x[2])|x[3])&x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[534] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[535] = ((((((x[3]&x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[536] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[537] = ((((((((x[1]|x[2])&x[3])&x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[538] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[539] = (((((((x[2]&x[3])&x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[540] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[541] = ((((((((x[1]&x[2])&x[3])&x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[542] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[543] = ((((x[5]|x[6])|x[7])|x[8])&x[9]);
assign y[544] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[545] = ((((((((x[1]|x[2])|x[3])|x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[546] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[547] = (((((((x[2]|x[3])|x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[548] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[549] = ((((((((x[1]&x[2])|x[3])|x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[550] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[551] = ((((((x[3]|x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[552] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[553] = ((((((((x[1]|x[2])&x[3])|x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[554] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[555] = (((((((x[2]&x[3])|x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[556] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[557] = ((((((((x[1]&x[2])&x[3])|x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[558] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[559] = (((((x[4]&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[560] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[561] = ((((((((x[1]|x[2])|x[3])&x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[562] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[563] = (((((((x[2]|x[3])&x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[564] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[565] = ((((((((x[1]&x[2])|x[3])&x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[566] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[567] = ((((((x[3]&x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[568] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[569] = ((((((((x[1]|x[2])&x[3])&x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[570] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[571] = (((((((x[2]&x[3])&x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[572] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[573] = ((((((((x[1]&x[2])&x[3])&x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[574] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])|x[6])|x[7])|x[8])&x[9]);
assign y[575] = (((x[6]|x[7])|x[8])&x[9]);
assign y[576] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[577] = ((((((((x[1]|x[2])|x[3])|x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[578] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[579] = (((((((x[2]|x[3])|x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[580] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[581] = ((((((((x[1]&x[2])|x[3])|x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[582] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[583] = ((((((x[3]|x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[584] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[585] = ((((((((x[1]|x[2])&x[3])|x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[586] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[587] = (((((((x[2]&x[3])|x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[588] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[589] = ((((((((x[1]&x[2])&x[3])|x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[590] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[591] = (((((x[4]|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[592] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[593] = ((((((((x[1]|x[2])|x[3])&x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[594] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[595] = (((((((x[2]|x[3])&x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[596] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[597] = ((((((((x[1]&x[2])|x[3])&x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[598] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[599] = ((((((x[3]&x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[600] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[601] = ((((((((x[1]|x[2])&x[3])&x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[602] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[603] = (((((((x[2]&x[3])&x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[604] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[605] = ((((((((x[1]&x[2])&x[3])&x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[606] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[607] = ((((x[5]&x[6])|x[7])|x[8])&x[9]);
assign y[608] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[609] = ((((((((x[1]|x[2])|x[3])|x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[610] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[611] = (((((((x[2]|x[3])|x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[612] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[613] = ((((((((x[1]&x[2])|x[3])|x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[614] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[615] = ((((((x[3]|x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[616] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[617] = ((((((((x[1]|x[2])&x[3])|x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[618] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[619] = (((((((x[2]&x[3])|x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[620] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[621] = ((((((((x[1]&x[2])&x[3])|x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[622] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[623] = (((((x[4]&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[624] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[625] = ((((((((x[1]|x[2])|x[3])&x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[626] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[627] = (((((((x[2]|x[3])&x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[628] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[629] = ((((((((x[1]&x[2])|x[3])&x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[630] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[631] = ((((((x[3]&x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[632] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[633] = ((((((((x[1]|x[2])&x[3])&x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[634] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[635] = (((((((x[2]&x[3])&x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[636] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[637] = ((((((((x[1]&x[2])&x[3])&x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[638] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])&x[6])|x[7])|x[8])&x[9]);
assign y[639] = ((x[7]|x[8])&x[9]);
assign y[640] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[641] = ((((((((x[1]|x[2])|x[3])|x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[642] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[643] = (((((((x[2]|x[3])|x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[644] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[645] = ((((((((x[1]&x[2])|x[3])|x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[646] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[647] = ((((((x[3]|x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[648] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[649] = ((((((((x[1]|x[2])&x[3])|x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[650] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[651] = (((((((x[2]&x[3])|x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[652] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[653] = ((((((((x[1]&x[2])&x[3])|x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[654] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[655] = (((((x[4]|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[656] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[657] = ((((((((x[1]|x[2])|x[3])&x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[658] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[659] = (((((((x[2]|x[3])&x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[660] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[661] = ((((((((x[1]&x[2])|x[3])&x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[662] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[663] = ((((((x[3]&x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[664] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[665] = ((((((((x[1]|x[2])&x[3])&x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[666] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[667] = (((((((x[2]&x[3])&x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[668] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[669] = ((((((((x[1]&x[2])&x[3])&x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[670] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[671] = ((((x[5]|x[6])&x[7])|x[8])&x[9]);
assign y[672] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[673] = ((((((((x[1]|x[2])|x[3])|x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[674] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[675] = (((((((x[2]|x[3])|x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[676] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[677] = ((((((((x[1]&x[2])|x[3])|x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[678] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[679] = ((((((x[3]|x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[680] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[681] = ((((((((x[1]|x[2])&x[3])|x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[682] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[683] = (((((((x[2]&x[3])|x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[684] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[685] = ((((((((x[1]&x[2])&x[3])|x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[686] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[687] = (((((x[4]&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[688] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[689] = ((((((((x[1]|x[2])|x[3])&x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[690] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[691] = (((((((x[2]|x[3])&x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[692] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[693] = ((((((((x[1]&x[2])|x[3])&x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[694] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[695] = ((((((x[3]&x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[696] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[697] = ((((((((x[1]|x[2])&x[3])&x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[698] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[699] = (((((((x[2]&x[3])&x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[700] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[701] = ((((((((x[1]&x[2])&x[3])&x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[702] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])|x[6])&x[7])|x[8])&x[9]);
assign y[703] = (((x[6]&x[7])|x[8])&x[9]);
assign y[704] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[705] = ((((((((x[1]|x[2])|x[3])|x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[706] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[707] = (((((((x[2]|x[3])|x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[708] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[709] = ((((((((x[1]&x[2])|x[3])|x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[710] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[711] = ((((((x[3]|x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[712] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[713] = ((((((((x[1]|x[2])&x[3])|x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[714] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[715] = (((((((x[2]&x[3])|x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[716] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[717] = ((((((((x[1]&x[2])&x[3])|x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[718] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[719] = (((((x[4]|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[720] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[721] = ((((((((x[1]|x[2])|x[3])&x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[722] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[723] = (((((((x[2]|x[3])&x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[724] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[725] = ((((((((x[1]&x[2])|x[3])&x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[726] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[727] = ((((((x[3]&x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[728] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[729] = ((((((((x[1]|x[2])&x[3])&x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[730] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[731] = (((((((x[2]&x[3])&x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[732] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[733] = ((((((((x[1]&x[2])&x[3])&x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[734] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[735] = ((((x[5]&x[6])&x[7])|x[8])&x[9]);
assign y[736] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[737] = ((((((((x[1]|x[2])|x[3])|x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[738] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[739] = (((((((x[2]|x[3])|x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[740] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[741] = ((((((((x[1]&x[2])|x[3])|x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[742] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[743] = ((((((x[3]|x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[744] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[745] = ((((((((x[1]|x[2])&x[3])|x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[746] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[747] = (((((((x[2]&x[3])|x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[748] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[749] = ((((((((x[1]&x[2])&x[3])|x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[750] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[751] = (((((x[4]&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[752] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[753] = ((((((((x[1]|x[2])|x[3])&x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[754] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[755] = (((((((x[2]|x[3])&x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[756] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[757] = ((((((((x[1]&x[2])|x[3])&x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[758] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[759] = ((((((x[3]&x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[760] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[761] = ((((((((x[1]|x[2])&x[3])&x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[762] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[763] = (((((((x[2]&x[3])&x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[764] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[765] = ((((((((x[1]&x[2])&x[3])&x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[766] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])&x[6])&x[7])|x[8])&x[9]);
assign y[767] = (x[8]&x[9]);
assign y[768] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[769] = ((((((((x[1]|x[2])|x[3])|x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[770] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[771] = (((((((x[2]|x[3])|x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[772] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[773] = ((((((((x[1]&x[2])|x[3])|x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[774] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[775] = ((((((x[3]|x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[776] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[777] = ((((((((x[1]|x[2])&x[3])|x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[778] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[779] = (((((((x[2]&x[3])|x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[780] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[781] = ((((((((x[1]&x[2])&x[3])|x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[782] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[783] = (((((x[4]|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[784] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[785] = ((((((((x[1]|x[2])|x[3])&x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[786] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[787] = (((((((x[2]|x[3])&x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[788] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[789] = ((((((((x[1]&x[2])|x[3])&x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[790] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[791] = ((((((x[3]&x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[792] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[793] = ((((((((x[1]|x[2])&x[3])&x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[794] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[795] = (((((((x[2]&x[3])&x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[796] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[797] = ((((((((x[1]&x[2])&x[3])&x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[798] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[799] = ((((x[5]|x[6])|x[7])&x[8])&x[9]);
assign y[800] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[801] = ((((((((x[1]|x[2])|x[3])|x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[802] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[803] = (((((((x[2]|x[3])|x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[804] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[805] = ((((((((x[1]&x[2])|x[3])|x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[806] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[807] = ((((((x[3]|x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[808] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[809] = ((((((((x[1]|x[2])&x[3])|x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[810] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[811] = (((((((x[2]&x[3])|x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[812] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[813] = ((((((((x[1]&x[2])&x[3])|x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[814] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[815] = (((((x[4]&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[816] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[817] = ((((((((x[1]|x[2])|x[3])&x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[818] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[819] = (((((((x[2]|x[3])&x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[820] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[821] = ((((((((x[1]&x[2])|x[3])&x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[822] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[823] = ((((((x[3]&x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[824] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[825] = ((((((((x[1]|x[2])&x[3])&x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[826] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[827] = (((((((x[2]&x[3])&x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[828] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[829] = ((((((((x[1]&x[2])&x[3])&x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[830] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])|x[6])|x[7])&x[8])&x[9]);
assign y[831] = (((x[6]|x[7])&x[8])&x[9]);
assign y[832] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[833] = ((((((((x[1]|x[2])|x[3])|x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[834] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[835] = (((((((x[2]|x[3])|x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[836] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[837] = ((((((((x[1]&x[2])|x[3])|x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[838] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[839] = ((((((x[3]|x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[840] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[841] = ((((((((x[1]|x[2])&x[3])|x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[842] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[843] = (((((((x[2]&x[3])|x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[844] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[845] = ((((((((x[1]&x[2])&x[3])|x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[846] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[847] = (((((x[4]|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[848] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[849] = ((((((((x[1]|x[2])|x[3])&x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[850] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[851] = (((((((x[2]|x[3])&x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[852] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[853] = ((((((((x[1]&x[2])|x[3])&x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[854] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[855] = ((((((x[3]&x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[856] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[857] = ((((((((x[1]|x[2])&x[3])&x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[858] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[859] = (((((((x[2]&x[3])&x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[860] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[861] = ((((((((x[1]&x[2])&x[3])&x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[862] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[863] = ((((x[5]&x[6])|x[7])&x[8])&x[9]);
assign y[864] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[865] = ((((((((x[1]|x[2])|x[3])|x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[866] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[867] = (((((((x[2]|x[3])|x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[868] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[869] = ((((((((x[1]&x[2])|x[3])|x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[870] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[871] = ((((((x[3]|x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[872] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[873] = ((((((((x[1]|x[2])&x[3])|x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[874] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[875] = (((((((x[2]&x[3])|x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[876] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[877] = ((((((((x[1]&x[2])&x[3])|x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[878] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[879] = (((((x[4]&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[880] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[881] = ((((((((x[1]|x[2])|x[3])&x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[882] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[883] = (((((((x[2]|x[3])&x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[884] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[885] = ((((((((x[1]&x[2])|x[3])&x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[886] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[887] = ((((((x[3]&x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[888] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[889] = ((((((((x[1]|x[2])&x[3])&x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[890] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[891] = (((((((x[2]&x[3])&x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[892] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[893] = ((((((((x[1]&x[2])&x[3])&x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[894] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])&x[6])|x[7])&x[8])&x[9]);
assign y[895] = ((x[7]&x[8])&x[9]);
assign y[896] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[897] = ((((((((x[1]|x[2])|x[3])|x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[898] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[899] = (((((((x[2]|x[3])|x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[900] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[901] = ((((((((x[1]&x[2])|x[3])|x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[902] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[903] = ((((((x[3]|x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[904] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[905] = ((((((((x[1]|x[2])&x[3])|x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[906] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[907] = (((((((x[2]&x[3])|x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[908] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[909] = ((((((((x[1]&x[2])&x[3])|x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[910] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[911] = (((((x[4]|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[912] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[913] = ((((((((x[1]|x[2])|x[3])&x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[914] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[915] = (((((((x[2]|x[3])&x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[916] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[917] = ((((((((x[1]&x[2])|x[3])&x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[918] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[919] = ((((((x[3]&x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[920] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[921] = ((((((((x[1]|x[2])&x[3])&x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[922] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[923] = (((((((x[2]&x[3])&x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[924] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[925] = ((((((((x[1]&x[2])&x[3])&x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[926] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[927] = ((((x[5]|x[6])&x[7])&x[8])&x[9]);
assign y[928] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[929] = ((((((((x[1]|x[2])|x[3])|x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[930] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[931] = (((((((x[2]|x[3])|x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[932] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[933] = ((((((((x[1]&x[2])|x[3])|x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[934] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[935] = ((((((x[3]|x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[936] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[937] = ((((((((x[1]|x[2])&x[3])|x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[938] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[939] = (((((((x[2]&x[3])|x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[940] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[941] = ((((((((x[1]&x[2])&x[3])|x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[942] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[943] = (((((x[4]&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[944] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[945] = ((((((((x[1]|x[2])|x[3])&x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[946] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[947] = (((((((x[2]|x[3])&x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[948] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[949] = ((((((((x[1]&x[2])|x[3])&x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[950] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[951] = ((((((x[3]&x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[952] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[953] = ((((((((x[1]|x[2])&x[3])&x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[954] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[955] = (((((((x[2]&x[3])&x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[956] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[957] = ((((((((x[1]&x[2])&x[3])&x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[958] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])|x[6])&x[7])&x[8])&x[9]);
assign y[959] = (((x[6]&x[7])&x[8])&x[9]);
assign y[960] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[961] = ((((((((x[1]|x[2])|x[3])|x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[962] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[963] = (((((((x[2]|x[3])|x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[964] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[965] = ((((((((x[1]&x[2])|x[3])|x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[966] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[967] = ((((((x[3]|x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[968] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[969] = ((((((((x[1]|x[2])&x[3])|x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[970] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[971] = (((((((x[2]&x[3])|x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[972] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[973] = ((((((((x[1]&x[2])&x[3])|x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[974] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[975] = (((((x[4]|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[976] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[977] = ((((((((x[1]|x[2])|x[3])&x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[978] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[979] = (((((((x[2]|x[3])&x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[980] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[981] = ((((((((x[1]&x[2])|x[3])&x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[982] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[983] = ((((((x[3]&x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[984] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[985] = ((((((((x[1]|x[2])&x[3])&x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[986] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[987] = (((((((x[2]&x[3])&x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[988] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[989] = ((((((((x[1]&x[2])&x[3])&x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[990] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])|x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[991] = ((((x[5]&x[6])&x[7])&x[8])&x[9]);
assign y[992] = (((((((((x[0]|x[1])|x[2])|x[3])|x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[993] = ((((((((x[1]|x[2])|x[3])|x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[994] = (((((((((x[0]&x[1])|x[2])|x[3])|x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[995] = (((((((x[2]|x[3])|x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[996] = (((((((((x[0]|x[1])&x[2])|x[3])|x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[997] = ((((((((x[1]&x[2])|x[3])|x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[998] = (((((((((x[0]&x[1])&x[2])|x[3])|x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[999] = ((((((x[3]|x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1000] = (((((((((x[0]|x[1])|x[2])&x[3])|x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1001] = ((((((((x[1]|x[2])&x[3])|x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1002] = (((((((((x[0]&x[1])|x[2])&x[3])|x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1003] = (((((((x[2]&x[3])|x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1004] = (((((((((x[0]|x[1])&x[2])&x[3])|x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1005] = ((((((((x[1]&x[2])&x[3])|x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1006] = (((((((((x[0]&x[1])&x[2])&x[3])|x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1007] = (((((x[4]&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1008] = (((((((((x[0]|x[1])|x[2])|x[3])&x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1009] = ((((((((x[1]|x[2])|x[3])&x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1010] = (((((((((x[0]&x[1])|x[2])|x[3])&x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1011] = (((((((x[2]|x[3])&x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1012] = (((((((((x[0]|x[1])&x[2])|x[3])&x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1013] = ((((((((x[1]&x[2])|x[3])&x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1014] = (((((((((x[0]&x[1])&x[2])|x[3])&x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1015] = ((((((x[3]&x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1016] = (((((((((x[0]|x[1])|x[2])&x[3])&x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1017] = ((((((((x[1]|x[2])&x[3])&x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1018] = (((((((((x[0]&x[1])|x[2])&x[3])&x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1019] = (((((((x[2]&x[3])&x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1020] = (((((((((x[0]|x[1])&x[2])&x[3])&x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1021] = ((((((((x[1]&x[2])&x[3])&x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1022] = (((((((((x[0]&x[1])&x[2])&x[3])&x[4])&x[5])&x[6])&x[7])&x[8])&x[9]);
assign y[1023] = 0;

endmodule 
